module gen_1Hz(input clk, input dcf_digital, output clk_1Hz);


